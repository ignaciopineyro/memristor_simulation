* MEMRISTOR CIRCUIT - MODEL pershin.sub

* DEPENDENCIES:
.include /home/ignaciopineyro/memristor_simulation/models/pershin.sub

* COMPONENTS:
V1 vin gnd sin 0 0.7 1   
xmem0 vin gnd l0 memristor

* ANALYSIS COMMANDS:
.tran 0.002 2 1e-09  uic

* CONTROL COMMANDS:
.control
run
set wr_vecnames
set wr_singlescale
wrdata /home/ignaciopineyro/memristor_simulation/simulation_results/pershin_simulations/di_francesco_vin_amplitude/vin_0.7.csv vin i(v1) l0
quit

.endc
.end
